VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_a51
  CLASS BLOCK ;
  FOREIGN wrapped_a51 ;
  ORIGIN 0.000 0.000 ;
  SIZE 380.000 BY 380.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.770 376.000 31.330 380.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 1.100 380.000 2.300 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 101.060 380.000 102.260 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 110.580 380.000 111.780 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 120.780 380.000 121.980 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 130.980 380.000 132.180 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 140.500 380.000 141.700 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 150.700 380.000 151.900 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 160.900 380.000 162.100 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 171.100 380.000 172.300 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 180.620 380.000 181.820 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 190.820 380.000 192.020 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 10.620 380.000 11.820 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 201.020 380.000 202.220 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 210.540 380.000 211.740 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 220.740 380.000 221.940 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 230.940 380.000 232.140 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 241.140 380.000 242.340 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 250.660 380.000 251.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 260.860 380.000 262.060 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 271.060 380.000 272.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 280.580 380.000 281.780 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 290.780 380.000 291.980 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 20.820 380.000 22.020 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 300.980 380.000 302.180 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 311.180 380.000 312.380 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 320.700 380.000 321.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 330.900 380.000 332.100 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 341.100 380.000 342.300 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 350.620 380.000 351.820 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 360.820 380.000 362.020 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 371.020 380.000 372.220 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 31.020 380.000 32.220 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 40.540 380.000 41.740 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 50.740 380.000 51.940 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 60.940 380.000 62.140 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 70.460 380.000 71.660 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 80.660 380.000 81.860 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 90.860 380.000 92.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 7.220 380.000 8.420 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 107.180 380.000 108.380 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 117.380 380.000 118.580 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 127.580 380.000 128.780 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 137.780 380.000 138.980 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 147.300 380.000 148.500 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 157.500 380.000 158.700 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 167.700 380.000 168.900 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 177.220 380.000 178.420 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 187.420 380.000 188.620 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 197.620 380.000 198.820 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 17.420 380.000 18.620 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 207.820 380.000 209.020 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 217.340 380.000 218.540 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 227.540 380.000 228.740 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 237.740 380.000 238.940 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 247.260 380.000 248.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 257.460 380.000 258.660 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 267.660 380.000 268.860 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 277.180 380.000 278.380 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 287.380 380.000 288.580 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 297.580 380.000 298.780 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 27.620 380.000 28.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 307.780 380.000 308.980 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 317.300 380.000 318.500 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 327.500 380.000 328.700 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 337.700 380.000 338.900 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 347.220 380.000 348.420 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 357.420 380.000 358.620 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 367.620 380.000 368.820 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 377.820 380.000 379.020 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 37.140 380.000 38.340 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 47.340 380.000 48.540 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 57.540 380.000 58.740 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 67.740 380.000 68.940 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 77.260 380.000 78.460 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 87.460 380.000 88.660 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 97.660 380.000 98.860 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 3.820 380.000 5.020 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 104.460 380.000 105.660 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 113.980 380.000 115.180 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 124.180 380.000 125.380 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 134.380 380.000 135.580 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 143.900 380.000 145.100 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 154.100 380.000 155.300 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 164.300 380.000 165.500 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 173.820 380.000 175.020 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 184.020 380.000 185.220 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 194.220 380.000 195.420 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 14.020 380.000 15.220 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 204.420 380.000 205.620 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 213.940 380.000 215.140 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 224.140 380.000 225.340 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 234.340 380.000 235.540 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 243.860 380.000 245.060 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 254.060 380.000 255.260 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 264.260 380.000 265.460 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 274.460 380.000 275.660 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 283.980 380.000 285.180 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 294.180 380.000 295.380 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 24.220 380.000 25.420 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 304.380 380.000 305.580 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 313.900 380.000 315.100 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 324.100 380.000 325.300 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 334.300 380.000 335.500 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 344.500 380.000 345.700 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 354.020 380.000 355.220 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 364.220 380.000 365.420 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 374.420 380.000 375.620 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 34.420 380.000 35.620 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 43.940 380.000 45.140 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 54.140 380.000 55.340 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 64.340 380.000 65.540 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 73.860 380.000 75.060 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 84.060 380.000 85.260 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 94.260 380.000 95.460 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.490 376.000 368.050 380.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.550 376.000 373.110 380.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 376.000 377.710 380.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 0.000 3.270 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.050 0.000 62.610 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 0.000 68.130 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 0.000 74.110 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 0.000 80.090 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.510 0.000 86.070 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.490 0.000 92.050 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 0.000 98.030 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.450 0.000 104.010 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 0.000 109.990 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 0.000 115.970 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 0.000 8.790 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 0.000 121.950 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.370 0.000 127.930 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.890 0.000 133.450 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.870 0.000 139.430 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 0.000 145.410 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.830 0.000 151.390 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.810 0.000 157.370 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.790 0.000 163.350 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.770 0.000 169.330 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 0.000 175.310 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 0.000 14.770 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.730 0.000 181.290 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 0.000 187.270 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 0.000 20.750 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 0.000 26.730 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 0.000 32.710 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 0.000 38.690 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 0.000 44.670 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.090 0.000 50.650 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 0.000 56.630 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 0.000 193.250 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.030 0.000 252.590 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.550 0.000 258.110 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.530 0.000 264.090 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.510 0.000 270.070 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.490 0.000 276.050 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.470 0.000 282.030 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.450 0.000 288.010 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.430 0.000 293.990 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.410 0.000 299.970 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.390 0.000 305.950 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.210 0.000 198.770 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.370 0.000 311.930 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.350 0.000 317.910 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.870 0.000 323.430 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.850 0.000 329.410 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.830 0.000 335.390 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.810 0.000 341.370 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.790 0.000 347.350 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.770 0.000 353.330 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.750 0.000 359.310 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 0.000 365.290 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.190 0.000 204.750 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.710 0.000 371.270 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.690 0.000 377.250 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.170 0.000 210.730 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.150 0.000 216.710 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.130 0.000 222.690 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.110 0.000 228.670 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.090 0.000 234.650 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.070 0.000 240.630 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.050 0.000 246.610 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.180 4.000 193.380 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.340 4.000 252.540 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.460 4.000 258.660 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.580 4.000 264.780 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.700 4.000 270.900 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.140 4.000 276.340 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.260 4.000 282.460 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.380 4.000 288.580 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.820 4.000 294.020 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.940 4.000 300.140 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.060 4.000 306.260 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.300 4.000 199.500 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.180 4.000 312.380 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.620 4.000 317.820 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.740 4.000 323.940 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.860 4.000 330.060 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.980 4.000 336.180 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.420 4.000 341.620 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.540 4.000 347.740 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.660 4.000 353.860 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.780 4.000 359.980 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.220 4.000 365.420 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.740 4.000 204.940 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.340 4.000 371.540 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.460 4.000 377.660 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.860 4.000 211.060 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.980 4.000 217.180 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.100 4.000 223.300 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.540 4.000 228.740 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.660 4.000 234.860 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.780 4.000 240.980 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.900 4.000 247.100 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.830 376.000 36.390 380.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 367.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 367.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 367.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 367.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 367.440 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.250 376.000 2.810 380.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.850 376.000 7.410 380.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 376.000 26.730 380.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.750 376.000 60.310 380.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.050 376.000 108.610 380.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 376.000 113.210 380.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.250 376.000 117.810 380.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 376.000 122.870 380.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.910 376.000 127.470 380.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 376.000 132.530 380.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.570 376.000 137.130 380.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 376.000 142.190 380.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.230 376.000 146.790 380.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 376.000 151.850 380.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 376.000 64.910 380.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.890 376.000 156.450 380.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.950 376.000 161.510 380.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.550 376.000 166.110 380.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.150 376.000 170.710 380.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.210 376.000 175.770 380.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 376.000 180.370 380.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.870 376.000 185.430 380.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.470 376.000 190.030 380.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.530 376.000 195.090 380.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.130 376.000 199.690 380.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.410 376.000 69.970 380.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.190 376.000 204.750 380.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.790 376.000 209.350 380.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 376.000 74.570 380.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 376.000 79.630 380.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 376.000 84.230 380.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.730 376.000 89.290 380.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.330 376.000 93.890 380.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.390 376.000 98.950 380.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 376.000 103.550 380.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.510 376.000 17.070 380.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.850 376.000 214.410 380.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.690 376.000 262.250 380.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.750 376.000 267.310 380.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.350 376.000 271.910 380.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.950 376.000 276.510 380.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.010 376.000 281.570 380.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.610 376.000 286.170 380.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.670 376.000 291.230 380.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.270 376.000 295.830 380.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.330 376.000 300.890 380.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.930 376.000 305.490 380.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.450 376.000 219.010 380.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 376.000 310.550 380.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.590 376.000 315.150 380.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.650 376.000 320.210 380.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.250 376.000 324.810 380.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.850 376.000 329.410 380.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.910 376.000 334.470 380.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.510 376.000 339.070 380.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.570 376.000 344.130 380.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.170 376.000 348.730 380.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.230 376.000 353.790 380.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.050 376.000 223.610 380.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.830 376.000 358.390 380.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 376.000 363.450 380.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.110 376.000 228.670 380.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.710 376.000 233.270 380.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.770 376.000 238.330 380.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.370 376.000 242.930 380.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.430 376.000 247.990 380.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.030 376.000 252.590 380.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.090 376.000 257.650 380.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.460 4.000 3.660 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.620 4.000 62.820 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.740 4.000 68.940 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.180 4.000 74.380 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.300 4.000 80.500 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.420 4.000 86.620 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.540 4.000 92.740 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.980 4.000 98.180 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.100 4.000 104.300 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.220 4.000 110.420 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.660 4.000 115.860 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.900 4.000 9.100 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.780 4.000 121.980 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.900 4.000 128.100 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.020 4.000 134.220 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.460 4.000 139.660 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.580 4.000 145.780 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.700 4.000 151.900 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.820 4.000 158.020 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.260 4.000 163.460 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.380 4.000 169.580 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.500 4.000 175.700 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.020 4.000 15.220 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.620 4.000 181.820 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.060 4.000 187.260 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.140 4.000 21.340 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.580 4.000 26.780 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.700 4.000 32.900 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.820 4.000 39.020 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.940 4.000 45.140 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.380 4.000 50.580 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.500 4.000 56.700 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 376.000 40.990 380.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.490 376.000 46.050 380.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.090 376.000 50.650 380.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.150 376.000 55.710 380.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.450 376.000 12.010 380.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.110 376.000 21.670 380.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 2.905 10.795 377.055 367.285 ;
      LAYER met1 ;
        RECT 0.070 6.500 377.590 376.340 ;
      LAYER met2 ;
        RECT 0.100 375.720 1.970 379.285 ;
        RECT 3.090 375.720 6.570 379.285 ;
        RECT 7.690 375.720 11.170 379.285 ;
        RECT 12.290 375.720 16.230 379.285 ;
        RECT 17.350 375.720 20.830 379.285 ;
        RECT 21.950 375.720 25.890 379.285 ;
        RECT 27.010 375.720 30.490 379.285 ;
        RECT 31.610 375.720 35.550 379.285 ;
        RECT 36.670 375.720 40.150 379.285 ;
        RECT 41.270 375.720 45.210 379.285 ;
        RECT 46.330 375.720 49.810 379.285 ;
        RECT 50.930 375.720 54.870 379.285 ;
        RECT 55.990 375.720 59.470 379.285 ;
        RECT 60.590 375.720 64.070 379.285 ;
        RECT 65.190 375.720 69.130 379.285 ;
        RECT 70.250 375.720 73.730 379.285 ;
        RECT 74.850 375.720 78.790 379.285 ;
        RECT 79.910 375.720 83.390 379.285 ;
        RECT 84.510 375.720 88.450 379.285 ;
        RECT 89.570 375.720 93.050 379.285 ;
        RECT 94.170 375.720 98.110 379.285 ;
        RECT 99.230 375.720 102.710 379.285 ;
        RECT 103.830 375.720 107.770 379.285 ;
        RECT 108.890 375.720 112.370 379.285 ;
        RECT 113.490 375.720 116.970 379.285 ;
        RECT 118.090 375.720 122.030 379.285 ;
        RECT 123.150 375.720 126.630 379.285 ;
        RECT 127.750 375.720 131.690 379.285 ;
        RECT 132.810 375.720 136.290 379.285 ;
        RECT 137.410 375.720 141.350 379.285 ;
        RECT 142.470 375.720 145.950 379.285 ;
        RECT 147.070 375.720 151.010 379.285 ;
        RECT 152.130 375.720 155.610 379.285 ;
        RECT 156.730 375.720 160.670 379.285 ;
        RECT 161.790 375.720 165.270 379.285 ;
        RECT 166.390 375.720 169.870 379.285 ;
        RECT 170.990 375.720 174.930 379.285 ;
        RECT 176.050 375.720 179.530 379.285 ;
        RECT 180.650 375.720 184.590 379.285 ;
        RECT 185.710 375.720 189.190 379.285 ;
        RECT 190.310 375.720 194.250 379.285 ;
        RECT 195.370 375.720 198.850 379.285 ;
        RECT 199.970 375.720 203.910 379.285 ;
        RECT 205.030 375.720 208.510 379.285 ;
        RECT 209.630 375.720 213.570 379.285 ;
        RECT 214.690 375.720 218.170 379.285 ;
        RECT 219.290 375.720 222.770 379.285 ;
        RECT 223.890 375.720 227.830 379.285 ;
        RECT 228.950 375.720 232.430 379.285 ;
        RECT 233.550 375.720 237.490 379.285 ;
        RECT 238.610 375.720 242.090 379.285 ;
        RECT 243.210 375.720 247.150 379.285 ;
        RECT 248.270 375.720 251.750 379.285 ;
        RECT 252.870 375.720 256.810 379.285 ;
        RECT 257.930 375.720 261.410 379.285 ;
        RECT 262.530 375.720 266.470 379.285 ;
        RECT 267.590 375.720 271.070 379.285 ;
        RECT 272.190 375.720 275.670 379.285 ;
        RECT 276.790 375.720 280.730 379.285 ;
        RECT 281.850 375.720 285.330 379.285 ;
        RECT 286.450 375.720 290.390 379.285 ;
        RECT 291.510 375.720 294.990 379.285 ;
        RECT 296.110 375.720 300.050 379.285 ;
        RECT 301.170 375.720 304.650 379.285 ;
        RECT 305.770 375.720 309.710 379.285 ;
        RECT 310.830 375.720 314.310 379.285 ;
        RECT 315.430 375.720 319.370 379.285 ;
        RECT 320.490 375.720 323.970 379.285 ;
        RECT 325.090 375.720 328.570 379.285 ;
        RECT 329.690 375.720 333.630 379.285 ;
        RECT 334.750 375.720 338.230 379.285 ;
        RECT 339.350 375.720 343.290 379.285 ;
        RECT 344.410 375.720 347.890 379.285 ;
        RECT 349.010 375.720 352.950 379.285 ;
        RECT 354.070 375.720 357.550 379.285 ;
        RECT 358.670 375.720 362.610 379.285 ;
        RECT 363.730 375.720 367.210 379.285 ;
        RECT 368.330 375.720 372.270 379.285 ;
        RECT 373.390 375.720 376.870 379.285 ;
        RECT 0.100 4.280 377.560 375.720 ;
        RECT 0.100 2.875 2.430 4.280 ;
        RECT 3.550 2.875 7.950 4.280 ;
        RECT 9.070 2.875 13.930 4.280 ;
        RECT 15.050 2.875 19.910 4.280 ;
        RECT 21.030 2.875 25.890 4.280 ;
        RECT 27.010 2.875 31.870 4.280 ;
        RECT 32.990 2.875 37.850 4.280 ;
        RECT 38.970 2.875 43.830 4.280 ;
        RECT 44.950 2.875 49.810 4.280 ;
        RECT 50.930 2.875 55.790 4.280 ;
        RECT 56.910 2.875 61.770 4.280 ;
        RECT 62.890 2.875 67.290 4.280 ;
        RECT 68.410 2.875 73.270 4.280 ;
        RECT 74.390 2.875 79.250 4.280 ;
        RECT 80.370 2.875 85.230 4.280 ;
        RECT 86.350 2.875 91.210 4.280 ;
        RECT 92.330 2.875 97.190 4.280 ;
        RECT 98.310 2.875 103.170 4.280 ;
        RECT 104.290 2.875 109.150 4.280 ;
        RECT 110.270 2.875 115.130 4.280 ;
        RECT 116.250 2.875 121.110 4.280 ;
        RECT 122.230 2.875 127.090 4.280 ;
        RECT 128.210 2.875 132.610 4.280 ;
        RECT 133.730 2.875 138.590 4.280 ;
        RECT 139.710 2.875 144.570 4.280 ;
        RECT 145.690 2.875 150.550 4.280 ;
        RECT 151.670 2.875 156.530 4.280 ;
        RECT 157.650 2.875 162.510 4.280 ;
        RECT 163.630 2.875 168.490 4.280 ;
        RECT 169.610 2.875 174.470 4.280 ;
        RECT 175.590 2.875 180.450 4.280 ;
        RECT 181.570 2.875 186.430 4.280 ;
        RECT 187.550 2.875 192.410 4.280 ;
        RECT 193.530 2.875 197.930 4.280 ;
        RECT 199.050 2.875 203.910 4.280 ;
        RECT 205.030 2.875 209.890 4.280 ;
        RECT 211.010 2.875 215.870 4.280 ;
        RECT 216.990 2.875 221.850 4.280 ;
        RECT 222.970 2.875 227.830 4.280 ;
        RECT 228.950 2.875 233.810 4.280 ;
        RECT 234.930 2.875 239.790 4.280 ;
        RECT 240.910 2.875 245.770 4.280 ;
        RECT 246.890 2.875 251.750 4.280 ;
        RECT 252.870 2.875 257.270 4.280 ;
        RECT 258.390 2.875 263.250 4.280 ;
        RECT 264.370 2.875 269.230 4.280 ;
        RECT 270.350 2.875 275.210 4.280 ;
        RECT 276.330 2.875 281.190 4.280 ;
        RECT 282.310 2.875 287.170 4.280 ;
        RECT 288.290 2.875 293.150 4.280 ;
        RECT 294.270 2.875 299.130 4.280 ;
        RECT 300.250 2.875 305.110 4.280 ;
        RECT 306.230 2.875 311.090 4.280 ;
        RECT 312.210 2.875 317.070 4.280 ;
        RECT 318.190 2.875 322.590 4.280 ;
        RECT 323.710 2.875 328.570 4.280 ;
        RECT 329.690 2.875 334.550 4.280 ;
        RECT 335.670 2.875 340.530 4.280 ;
        RECT 341.650 2.875 346.510 4.280 ;
        RECT 347.630 2.875 352.490 4.280 ;
        RECT 353.610 2.875 358.470 4.280 ;
        RECT 359.590 2.875 364.450 4.280 ;
        RECT 365.570 2.875 370.430 4.280 ;
        RECT 371.550 2.875 376.410 4.280 ;
        RECT 377.530 2.875 377.560 4.280 ;
      LAYER met3 ;
        RECT 0.270 378.060 375.600 379.265 ;
        RECT 4.400 377.420 375.600 378.060 ;
        RECT 4.400 376.060 376.000 377.420 ;
        RECT 0.270 376.020 376.000 376.060 ;
        RECT 0.270 374.020 375.600 376.020 ;
        RECT 0.270 372.620 376.000 374.020 ;
        RECT 0.270 371.940 375.600 372.620 ;
        RECT 4.400 370.620 375.600 371.940 ;
        RECT 4.400 369.940 376.000 370.620 ;
        RECT 0.270 369.220 376.000 369.940 ;
        RECT 0.270 367.220 375.600 369.220 ;
        RECT 0.270 365.820 376.000 367.220 ;
        RECT 4.400 363.820 375.600 365.820 ;
        RECT 0.270 362.420 376.000 363.820 ;
        RECT 0.270 360.420 375.600 362.420 ;
        RECT 0.270 360.380 376.000 360.420 ;
        RECT 4.400 359.020 376.000 360.380 ;
        RECT 4.400 358.380 375.600 359.020 ;
        RECT 0.270 357.020 375.600 358.380 ;
        RECT 0.270 355.620 376.000 357.020 ;
        RECT 0.270 354.260 375.600 355.620 ;
        RECT 4.400 353.620 375.600 354.260 ;
        RECT 4.400 352.260 376.000 353.620 ;
        RECT 0.270 352.220 376.000 352.260 ;
        RECT 0.270 350.220 375.600 352.220 ;
        RECT 0.270 348.820 376.000 350.220 ;
        RECT 0.270 348.140 375.600 348.820 ;
        RECT 4.400 346.820 375.600 348.140 ;
        RECT 4.400 346.140 376.000 346.820 ;
        RECT 0.270 346.100 376.000 346.140 ;
        RECT 0.270 344.100 375.600 346.100 ;
        RECT 0.270 342.700 376.000 344.100 ;
        RECT 0.270 342.020 375.600 342.700 ;
        RECT 4.400 340.700 375.600 342.020 ;
        RECT 4.400 340.020 376.000 340.700 ;
        RECT 0.270 339.300 376.000 340.020 ;
        RECT 0.270 337.300 375.600 339.300 ;
        RECT 0.270 336.580 376.000 337.300 ;
        RECT 4.400 335.900 376.000 336.580 ;
        RECT 4.400 334.580 375.600 335.900 ;
        RECT 0.270 333.900 375.600 334.580 ;
        RECT 0.270 332.500 376.000 333.900 ;
        RECT 0.270 330.500 375.600 332.500 ;
        RECT 0.270 330.460 376.000 330.500 ;
        RECT 4.400 329.100 376.000 330.460 ;
        RECT 4.400 328.460 375.600 329.100 ;
        RECT 0.270 327.100 375.600 328.460 ;
        RECT 0.270 325.700 376.000 327.100 ;
        RECT 0.270 324.340 375.600 325.700 ;
        RECT 4.400 323.700 375.600 324.340 ;
        RECT 4.400 322.340 376.000 323.700 ;
        RECT 0.270 322.300 376.000 322.340 ;
        RECT 0.270 320.300 375.600 322.300 ;
        RECT 0.270 318.900 376.000 320.300 ;
        RECT 0.270 318.220 375.600 318.900 ;
        RECT 4.400 316.900 375.600 318.220 ;
        RECT 4.400 316.220 376.000 316.900 ;
        RECT 0.270 315.500 376.000 316.220 ;
        RECT 0.270 313.500 375.600 315.500 ;
        RECT 0.270 312.780 376.000 313.500 ;
        RECT 4.400 310.780 375.600 312.780 ;
        RECT 0.270 309.380 376.000 310.780 ;
        RECT 0.270 307.380 375.600 309.380 ;
        RECT 0.270 306.660 376.000 307.380 ;
        RECT 4.400 305.980 376.000 306.660 ;
        RECT 4.400 304.660 375.600 305.980 ;
        RECT 0.270 303.980 375.600 304.660 ;
        RECT 0.270 302.580 376.000 303.980 ;
        RECT 0.270 300.580 375.600 302.580 ;
        RECT 0.270 300.540 376.000 300.580 ;
        RECT 4.400 299.180 376.000 300.540 ;
        RECT 4.400 298.540 375.600 299.180 ;
        RECT 0.270 297.180 375.600 298.540 ;
        RECT 0.270 295.780 376.000 297.180 ;
        RECT 0.270 294.420 375.600 295.780 ;
        RECT 4.400 293.780 375.600 294.420 ;
        RECT 4.400 292.420 376.000 293.780 ;
        RECT 0.270 292.380 376.000 292.420 ;
        RECT 0.270 290.380 375.600 292.380 ;
        RECT 0.270 288.980 376.000 290.380 ;
        RECT 4.400 286.980 375.600 288.980 ;
        RECT 0.270 285.580 376.000 286.980 ;
        RECT 0.270 283.580 375.600 285.580 ;
        RECT 0.270 282.860 376.000 283.580 ;
        RECT 4.400 282.180 376.000 282.860 ;
        RECT 4.400 280.860 375.600 282.180 ;
        RECT 0.270 280.180 375.600 280.860 ;
        RECT 0.270 278.780 376.000 280.180 ;
        RECT 0.270 276.780 375.600 278.780 ;
        RECT 0.270 276.740 376.000 276.780 ;
        RECT 4.400 276.060 376.000 276.740 ;
        RECT 4.400 274.740 375.600 276.060 ;
        RECT 0.270 274.060 375.600 274.740 ;
        RECT 0.270 272.660 376.000 274.060 ;
        RECT 0.270 271.300 375.600 272.660 ;
        RECT 4.400 270.660 375.600 271.300 ;
        RECT 4.400 269.300 376.000 270.660 ;
        RECT 0.270 269.260 376.000 269.300 ;
        RECT 0.270 267.260 375.600 269.260 ;
        RECT 0.270 265.860 376.000 267.260 ;
        RECT 0.270 265.180 375.600 265.860 ;
        RECT 4.400 263.860 375.600 265.180 ;
        RECT 4.400 263.180 376.000 263.860 ;
        RECT 0.270 262.460 376.000 263.180 ;
        RECT 0.270 260.460 375.600 262.460 ;
        RECT 0.270 259.060 376.000 260.460 ;
        RECT 4.400 257.060 375.600 259.060 ;
        RECT 0.270 255.660 376.000 257.060 ;
        RECT 0.270 253.660 375.600 255.660 ;
        RECT 0.270 252.940 376.000 253.660 ;
        RECT 4.400 252.260 376.000 252.940 ;
        RECT 4.400 250.940 375.600 252.260 ;
        RECT 0.270 250.260 375.600 250.940 ;
        RECT 0.270 248.860 376.000 250.260 ;
        RECT 0.270 247.500 375.600 248.860 ;
        RECT 4.400 246.860 375.600 247.500 ;
        RECT 4.400 245.500 376.000 246.860 ;
        RECT 0.270 245.460 376.000 245.500 ;
        RECT 0.270 243.460 375.600 245.460 ;
        RECT 0.270 242.740 376.000 243.460 ;
        RECT 0.270 241.380 375.600 242.740 ;
        RECT 4.400 240.740 375.600 241.380 ;
        RECT 4.400 239.380 376.000 240.740 ;
        RECT 0.270 239.340 376.000 239.380 ;
        RECT 0.270 237.340 375.600 239.340 ;
        RECT 0.270 235.940 376.000 237.340 ;
        RECT 0.270 235.260 375.600 235.940 ;
        RECT 4.400 233.940 375.600 235.260 ;
        RECT 4.400 233.260 376.000 233.940 ;
        RECT 0.270 232.540 376.000 233.260 ;
        RECT 0.270 230.540 375.600 232.540 ;
        RECT 0.270 229.140 376.000 230.540 ;
        RECT 4.400 227.140 375.600 229.140 ;
        RECT 0.270 225.740 376.000 227.140 ;
        RECT 0.270 223.740 375.600 225.740 ;
        RECT 0.270 223.700 376.000 223.740 ;
        RECT 4.400 222.340 376.000 223.700 ;
        RECT 4.400 221.700 375.600 222.340 ;
        RECT 0.270 220.340 375.600 221.700 ;
        RECT 0.270 218.940 376.000 220.340 ;
        RECT 0.270 217.580 375.600 218.940 ;
        RECT 4.400 216.940 375.600 217.580 ;
        RECT 4.400 215.580 376.000 216.940 ;
        RECT 0.270 215.540 376.000 215.580 ;
        RECT 0.270 213.540 375.600 215.540 ;
        RECT 0.270 212.140 376.000 213.540 ;
        RECT 0.270 211.460 375.600 212.140 ;
        RECT 4.400 210.140 375.600 211.460 ;
        RECT 4.400 209.460 376.000 210.140 ;
        RECT 0.270 209.420 376.000 209.460 ;
        RECT 0.270 207.420 375.600 209.420 ;
        RECT 0.270 206.020 376.000 207.420 ;
        RECT 0.270 205.340 375.600 206.020 ;
        RECT 4.400 204.020 375.600 205.340 ;
        RECT 4.400 203.340 376.000 204.020 ;
        RECT 0.270 202.620 376.000 203.340 ;
        RECT 0.270 200.620 375.600 202.620 ;
        RECT 0.270 199.900 376.000 200.620 ;
        RECT 4.400 199.220 376.000 199.900 ;
        RECT 4.400 197.900 375.600 199.220 ;
        RECT 0.270 197.220 375.600 197.900 ;
        RECT 0.270 195.820 376.000 197.220 ;
        RECT 0.270 193.820 375.600 195.820 ;
        RECT 0.270 193.780 376.000 193.820 ;
        RECT 4.400 192.420 376.000 193.780 ;
        RECT 4.400 191.780 375.600 192.420 ;
        RECT 0.270 190.420 375.600 191.780 ;
        RECT 0.270 189.020 376.000 190.420 ;
        RECT 0.270 187.660 375.600 189.020 ;
        RECT 4.400 187.020 375.600 187.660 ;
        RECT 4.400 185.660 376.000 187.020 ;
        RECT 0.270 185.620 376.000 185.660 ;
        RECT 0.270 183.620 375.600 185.620 ;
        RECT 0.270 182.220 376.000 183.620 ;
        RECT 4.400 180.220 375.600 182.220 ;
        RECT 0.270 178.820 376.000 180.220 ;
        RECT 0.270 176.820 375.600 178.820 ;
        RECT 0.270 176.100 376.000 176.820 ;
        RECT 4.400 175.420 376.000 176.100 ;
        RECT 4.400 174.100 375.600 175.420 ;
        RECT 0.270 173.420 375.600 174.100 ;
        RECT 0.270 172.700 376.000 173.420 ;
        RECT 0.270 170.700 375.600 172.700 ;
        RECT 0.270 169.980 376.000 170.700 ;
        RECT 4.400 169.300 376.000 169.980 ;
        RECT 4.400 167.980 375.600 169.300 ;
        RECT 0.270 167.300 375.600 167.980 ;
        RECT 0.270 165.900 376.000 167.300 ;
        RECT 0.270 163.900 375.600 165.900 ;
        RECT 0.270 163.860 376.000 163.900 ;
        RECT 4.400 162.500 376.000 163.860 ;
        RECT 4.400 161.860 375.600 162.500 ;
        RECT 0.270 160.500 375.600 161.860 ;
        RECT 0.270 159.100 376.000 160.500 ;
        RECT 0.270 158.420 375.600 159.100 ;
        RECT 4.400 157.100 375.600 158.420 ;
        RECT 4.400 156.420 376.000 157.100 ;
        RECT 0.270 155.700 376.000 156.420 ;
        RECT 0.270 153.700 375.600 155.700 ;
        RECT 0.270 152.300 376.000 153.700 ;
        RECT 4.400 150.300 375.600 152.300 ;
        RECT 0.270 148.900 376.000 150.300 ;
        RECT 0.270 146.900 375.600 148.900 ;
        RECT 0.270 146.180 376.000 146.900 ;
        RECT 4.400 145.500 376.000 146.180 ;
        RECT 4.400 144.180 375.600 145.500 ;
        RECT 0.270 143.500 375.600 144.180 ;
        RECT 0.270 142.100 376.000 143.500 ;
        RECT 0.270 140.100 375.600 142.100 ;
        RECT 0.270 140.060 376.000 140.100 ;
        RECT 4.400 139.380 376.000 140.060 ;
        RECT 4.400 138.060 375.600 139.380 ;
        RECT 0.270 137.380 375.600 138.060 ;
        RECT 0.270 135.980 376.000 137.380 ;
        RECT 0.270 134.620 375.600 135.980 ;
        RECT 4.400 133.980 375.600 134.620 ;
        RECT 4.400 132.620 376.000 133.980 ;
        RECT 0.270 132.580 376.000 132.620 ;
        RECT 0.270 130.580 375.600 132.580 ;
        RECT 0.270 129.180 376.000 130.580 ;
        RECT 0.270 128.500 375.600 129.180 ;
        RECT 4.400 127.180 375.600 128.500 ;
        RECT 4.400 126.500 376.000 127.180 ;
        RECT 0.270 125.780 376.000 126.500 ;
        RECT 0.270 123.780 375.600 125.780 ;
        RECT 0.270 122.380 376.000 123.780 ;
        RECT 4.400 120.380 375.600 122.380 ;
        RECT 0.270 118.980 376.000 120.380 ;
        RECT 0.270 116.980 375.600 118.980 ;
        RECT 0.270 116.260 376.000 116.980 ;
        RECT 4.400 115.580 376.000 116.260 ;
        RECT 4.400 114.260 375.600 115.580 ;
        RECT 0.270 113.580 375.600 114.260 ;
        RECT 0.270 112.180 376.000 113.580 ;
        RECT 0.270 110.820 375.600 112.180 ;
        RECT 4.400 110.180 375.600 110.820 ;
        RECT 4.400 108.820 376.000 110.180 ;
        RECT 0.270 108.780 376.000 108.820 ;
        RECT 0.270 106.780 375.600 108.780 ;
        RECT 0.270 106.060 376.000 106.780 ;
        RECT 0.270 104.700 375.600 106.060 ;
        RECT 4.400 104.060 375.600 104.700 ;
        RECT 4.400 102.700 376.000 104.060 ;
        RECT 0.270 102.660 376.000 102.700 ;
        RECT 0.270 100.660 375.600 102.660 ;
        RECT 0.270 99.260 376.000 100.660 ;
        RECT 0.270 98.580 375.600 99.260 ;
        RECT 4.400 97.260 375.600 98.580 ;
        RECT 4.400 96.580 376.000 97.260 ;
        RECT 0.270 95.860 376.000 96.580 ;
        RECT 0.270 93.860 375.600 95.860 ;
        RECT 0.270 93.140 376.000 93.860 ;
        RECT 4.400 92.460 376.000 93.140 ;
        RECT 4.400 91.140 375.600 92.460 ;
        RECT 0.270 90.460 375.600 91.140 ;
        RECT 0.270 89.060 376.000 90.460 ;
        RECT 0.270 87.060 375.600 89.060 ;
        RECT 0.270 87.020 376.000 87.060 ;
        RECT 4.400 85.660 376.000 87.020 ;
        RECT 4.400 85.020 375.600 85.660 ;
        RECT 0.270 83.660 375.600 85.020 ;
        RECT 0.270 82.260 376.000 83.660 ;
        RECT 0.270 80.900 375.600 82.260 ;
        RECT 4.400 80.260 375.600 80.900 ;
        RECT 4.400 78.900 376.000 80.260 ;
        RECT 0.270 78.860 376.000 78.900 ;
        RECT 0.270 76.860 375.600 78.860 ;
        RECT 0.270 75.460 376.000 76.860 ;
        RECT 0.270 74.780 375.600 75.460 ;
        RECT 4.400 73.460 375.600 74.780 ;
        RECT 4.400 72.780 376.000 73.460 ;
        RECT 0.270 72.060 376.000 72.780 ;
        RECT 0.270 70.060 375.600 72.060 ;
        RECT 0.270 69.340 376.000 70.060 ;
        RECT 4.400 67.340 375.600 69.340 ;
        RECT 0.270 65.940 376.000 67.340 ;
        RECT 0.270 63.940 375.600 65.940 ;
        RECT 0.270 63.220 376.000 63.940 ;
        RECT 4.400 62.540 376.000 63.220 ;
        RECT 4.400 61.220 375.600 62.540 ;
        RECT 0.270 60.540 375.600 61.220 ;
        RECT 0.270 59.140 376.000 60.540 ;
        RECT 0.270 57.140 375.600 59.140 ;
        RECT 0.270 57.100 376.000 57.140 ;
        RECT 4.400 55.740 376.000 57.100 ;
        RECT 4.400 55.100 375.600 55.740 ;
        RECT 0.270 53.740 375.600 55.100 ;
        RECT 0.270 52.340 376.000 53.740 ;
        RECT 0.270 50.980 375.600 52.340 ;
        RECT 4.400 50.340 375.600 50.980 ;
        RECT 4.400 48.980 376.000 50.340 ;
        RECT 0.270 48.940 376.000 48.980 ;
        RECT 0.270 46.940 375.600 48.940 ;
        RECT 0.270 45.540 376.000 46.940 ;
        RECT 4.400 43.540 375.600 45.540 ;
        RECT 0.270 42.140 376.000 43.540 ;
        RECT 0.270 40.140 375.600 42.140 ;
        RECT 0.270 39.420 376.000 40.140 ;
        RECT 4.400 38.740 376.000 39.420 ;
        RECT 4.400 37.420 375.600 38.740 ;
        RECT 0.270 36.740 375.600 37.420 ;
        RECT 0.270 36.020 376.000 36.740 ;
        RECT 0.270 34.020 375.600 36.020 ;
        RECT 0.270 33.300 376.000 34.020 ;
        RECT 4.400 32.620 376.000 33.300 ;
        RECT 4.400 31.300 375.600 32.620 ;
        RECT 0.270 30.620 375.600 31.300 ;
        RECT 0.270 29.220 376.000 30.620 ;
        RECT 0.270 27.220 375.600 29.220 ;
        RECT 0.270 27.180 376.000 27.220 ;
        RECT 4.400 25.820 376.000 27.180 ;
        RECT 4.400 25.180 375.600 25.820 ;
        RECT 0.270 23.820 375.600 25.180 ;
        RECT 0.270 22.420 376.000 23.820 ;
        RECT 0.270 21.740 375.600 22.420 ;
        RECT 4.400 20.420 375.600 21.740 ;
        RECT 4.400 19.740 376.000 20.420 ;
        RECT 0.270 19.020 376.000 19.740 ;
        RECT 0.270 17.020 375.600 19.020 ;
        RECT 0.270 15.620 376.000 17.020 ;
        RECT 4.400 13.620 375.600 15.620 ;
        RECT 0.270 12.220 376.000 13.620 ;
        RECT 0.270 10.220 375.600 12.220 ;
        RECT 0.270 9.500 376.000 10.220 ;
        RECT 4.400 8.820 376.000 9.500 ;
        RECT 4.400 7.500 375.600 8.820 ;
        RECT 0.270 6.820 375.600 7.500 ;
        RECT 0.270 5.420 376.000 6.820 ;
        RECT 0.270 4.060 375.600 5.420 ;
        RECT 4.400 3.420 375.600 4.060 ;
        RECT 4.400 2.895 376.000 3.420 ;
      LAYER met4 ;
        RECT 0.295 367.840 279.385 379.265 ;
        RECT 0.295 11.055 20.640 367.840 ;
        RECT 23.040 11.055 97.440 367.840 ;
        RECT 99.840 11.055 174.240 367.840 ;
        RECT 176.640 11.055 251.040 367.840 ;
        RECT 253.440 11.055 279.385 367.840 ;
  END
END wrapped_a51
END LIBRARY

